//-----------------------------------------------------------------------------
// Testbench
//
// This testbench sets up and runs a simulation of the single-cycle RV32I CPU.
// It generates the system clock and reset signal, instantiates the top-level
// processor module, and runs a loaded RISC-V program from memory. The testbench
// is used to verify correct instruction execution, data movement, and overall
// CPU behavior over multiple cycles.
//
// File Contributor(s): 
//-----------------------------------------------------------------------------
