//-----------------------------------------------------------------------------
// Top Level Module
//
// This module instantiates and connects all core components of a single-cycle
// 32-bit RV32I RISC-V processor, including the program counter, instruction
// decoder, register file, ALU, control units, and memory interface.
//
// File Contributor(s):
//-----------------------------------------------------------------------------
